lpm_add_sub0_inst : lpm_add_sub0 PORT MAP (
		datab	 => datab_sig,
		result	 => result_sig
	);
