altaccumulate2_inst : altaccumulate2 PORT MAP (
		aclr	 => aclr_sig,
		clken	 => clken_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		result	 => result_sig
	);
