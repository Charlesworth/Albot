altaccumulate0_inst : altaccumulate0 PORT MAP (
		aclr	 => aclr_sig,
		clken	 => clken_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		cout	 => cout_sig,
		result	 => result_sig
	);
