lpm_compare2_inst : lpm_compare2 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		AgeB	 => AgeB_sig
	);
