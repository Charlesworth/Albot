lpm_add_sub1_inst : lpm_add_sub1 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		cout	 => cout_sig,
		result	 => result_sig
	);
