--*****************************************
-- (c) Phil Culverhouse, 2006
--
-- All rights reserved
-- 
-- CHANGES: 
-- 30.06.07 increased CoulumnCounter to 11 bits to avoid overflo during row
-- 30.06.07 added Hsync to AccumulateSignal to avoid accumulating pixels outside of Href
-- 02.07.07  fixed bug in YUV state machine allocated wrong timing to pixel enables
--
--********************************************

LIBRARY ieee;
USE ieee.std_logic_1164.all;
-- not both this and below -- USE ieee.std_logic_arith.all;
--use IEEE.numeric_bit.all; -- for integer to bit_vector conversion
use IEEE.numeric_std.all; -- for integer to bit_vector conversion

-- VGA std format 640 by 480 pixels in a frame
-- register them, count line by line
-- 

ENTITY SyncProcessor IS
	PORT
	(
		Clk 		 : IN  std_logic;
		Vsync 		 : IN std_logic;
		Hsync		 : IN std_logic;
		TrainFlag 	 : IN  std_logic; -- from debounced user switch input
		Aclr		 : IN std_logic; -- hold decode of pixel colour 01==red, 10==green, 11==blue
		YUV			 : out unsigned (2 downto 0); -- values R, G and B 4 pixels in a stream 000 is only set during Vsync
		Row			 : out unsigned (8 downto 0); -- 480 == 256+128+64 ie. "111100000"
		Column		 : out unsigned (10 downto 0); -- 640 == 512+128 ie. "1010000000"
		AccumulateSIGNAL : out std_logic; -- is HIGH during hysnc's within a frame, reset by Vsync
		CalculateSIGNAL : out std_logic; -- is HIGH during gap between last hysnc in a frame, reset by Vsync
		FirstROW	: out std_logic; -- true for first row in frame
		LastROW		: out std_logic; -- true for last row in frame
		WindowROW	: out std_logic; -- true for valid ROWs in specified processing window
		WindowCOLUMN: out std_logic;  -- true for valid COLUMNs in specified processing window
		TrainFLAGsynced:out std_logic; -- the user input TrainFLAG now sync'd to one frame only
		YUVclk: out std_logic;
		Yclk: out std_logic;
		Uclk: out std_logic;
		Y1clk: out std_logic;
		Vclk: out std_logic -- BGRG pixel seq.
		
	);
END SyncProcessor;


-- first register the pixel stream
ARCHITECTURE SyncProcessor_v1 OF SyncProcessor IS

	constant VGAmaxROW: natural := 480;
	constant VGAmaxCOLUMN: natural := 640*2; -- 1280 pixels in a line (UY for pixel N and then VY for pixel N+1)
	
	--##########################################################################################
	-- processing window size
	constant RwinSTARTc: natural	:= (VGAmaxROW/2)-3; -- was -50; -- for inverted connector, but upright camera --(240-25);
	constant RwinENDc: natural	:= (VGAmaxROW/2)+3; --(240+25);
	constant CwinSTARTc: natural	:= ((VGAmaxCOLUMN/2)-12);-- centre of FOV
	constant CwinENDc: natural	:= ((VGAmaxCOLUMN/2)+12); 
	
	--##########################################################################################	
	shared variable FrameCounter: natural :=0; -- counts frames up to limit of integer range
	signal YUV_Cstate, YUV_Nstate: unsigned (2 downto 0); -- natural range 0 to 3; -- was unsigned (2 downto 0); 
	signal RowCounter : natural range 0 to VGAmaxROW; --was unsigned (8 downto 0);
	signal ColumnCounter: natural range 0 to VGAmaxCOLUMN; -- was unsigned (9 downto 0);
	signal LastROWint:  std_logic; -- true for last row in frame
	signal RowCENTRE,ColumnCENTRE: std_logic;
	signal INFrameFLAGint: std_logic; -- '1' for all Hsync rows in a frame
	signal CalculateSIGNALint: std_logic; 
	signal STOP: std_logic :='1'; -- used to enable the counter, hence cleared to stop it.
	signal TrainFLAGstart,resetFLAG: std_logic; -- sync's start of training with Vsync 
	signal TrainDELAYED, TrainDELAYEDmore: std_logic;
	
	component dff port(d,clk,clrn,prn:in std_logic; q:out std_logic);end component;


BEGIN
	Row <= to_unsigned(Rowcounter,9); -- was RowCounter ; -- WAS (to_unsigned(Rowcounter,9)); -- convert integer to bit_vector!
	---PC 30.06.07  Column <= to_unsigned(Columncounter,10); -- was ColumnCounter; -- was (to_unsigned(Columncounter,10));
	Column <= to_unsigned(Columncounter,11); -- was ColumnCounter; -- was (to_unsigned(Columncounter,10));
	YUV <= YUV_Cstate; -- was to_unsigned(YUVcounter,3); --- was YUVcounter; 
	LastROW <= LastROWint and Hsync; -- ensure it does not stay true until next Vsync.
	
	
	
	-- now the sequencer for generating the syncronised TrainFLAG to ensure TrainFLAG only lasts one frame
u1: dff port map('1',TrainFLAG,not(STOP),'1',TrainDELAYED);-- train for one frame only
u2: dff port map(TrainDELAYED,Vsync, not(STOP),'1',TrainDELAYEDmore);-- train for one frame only
u3: dff port map(TrainDELAYEDmore,Vsync, '1','1',STOP);-- train for one frame only
	TrainFLAGsynced <= TrainDELAYEDmore; -- debug 
	--PC 30.06.07 AccumulateSIGNAL <=  INFrameFLAGint and not(Vsync) and (not(CalculateSIGNALint)); -- (not(LastROWint and INFrameFLAGint)); -- ensure it does not stay true until next Vsync.
	AccumulateSIGNAL <=  INFrameFLAGint and not(Vsync) and (not(CalculateSIGNALint)) and Hsync; -- (not(LastROWint and INFrameFLAGint)); -- ensure it does not stay true until next Vsync.
u4: dff port map('1',LastROWint, INFrameFLAGint,'1',CalculateSIGNALint);-- train for one frame only
	CalculateSIGNAL <= CalculateSIGNALint; -- LastROWint and INFrameFLAGint; -- ensure it does not stay true until next Vsync.

	-- sequential processes belowand Hsync; -- (not(LastROWint and INFrameFLAGint)); -- 
	---------------------------------------------------------------------------
	SYNC: PROCESS (Clk, Hsync)
	BEGIN
		if 	(Clk'event) and (Clk = '1')  then -- PC 04.08.06 was '1'
			if (Hsync = '1') then
				ColumnCounter <= ColumnCounter + 1;
	     	elsif (Hsync = '0')then
				ColumnCounter <= 0; 
			end if;
		end if;
	END PROCESS SYNC ;
	---------------------------------------------------------------------------
	HsyncCOUNT: process (Hsync, Vsync, Rowcounter)
	begin
		if  (Hsync'event) and (Hsync = '1') then -- increment row counter every line 
			RowCounter <= RowCounter +1;
			INframeFLAGint <= '1';
			if RowCounter > VGAmaxROW then
				RowCounter <= 0;
				end if;			
		end if;
		if (Vsync = '1') then
		    RowCounter <= 0; --"000000000";
			INframeFLAGint <= '0';
			FirstROW <= '0';
			LastROWint <= '0';
		end if;
		case RowCounter is
			when 1 =>
				FirstROW <= '1';
				LastROWint <= '0';
			when VGAmaxROW =>
				FirstROW <= '0';
				LastROWint <= '1';
			when others =>
				FirstROW <= '0';
				LastROWint <= '0';
			end case;
	end process HsyncCOUNT;
	---------------------------------------------------------------------------
	VsyncCOUNT: process (Vsync)
	begin
		if  (Vsync'event) and (Vsync = '1') then -- increment row counter every line 
			Framecounter := Framecounter +1;
		end if;
	end process VsyncCOUNT;
	---------------------------------------------------------------------------
	-- used to output a centre of frame pulse FOR TRAINING
	RowPULSE: process (RowCounter, Hsync)
	begin
		if (RowCounter >= RwinSTARTc)and (RowCounter <= RwinENDc) then --and (Hsync= '1') then --240
			WindowROW <= '1';
		else 
			WindowROW <= '0';
		end if;
	end process RowPULSE;	
	---------------------------------------------------------------------------
	ColumnPULSE: process (ColumnCounter, Hsync)
	begin
		if (ColumnCounter >= CwinSTARTc) and (ColumnCounter <= CwinENDc) then -- was and (Hsync = '1') then --1
			WindowCOLUMN <= '1';
		else 
			WindowCOLUMN <= '0';
		end if;
	end process ColumnPULSE;
	---------------------------------------------------------------------------
		---------------------------------------------------------------------------
	YUVCLOCK: process (clk, Hsync, YUV_Nstate) -- clk pixels on 4th pixel, so they are stable for 4 pixel clks.
	begin
		if (Hsync='0') then
			YUV_Cstate <="000";
		elsif (clk'event) and (clk = '1') then -- PC 03.07.07 was '0', as pixels change on falling edge, but FSM must change with regstered pixels
			YUV_Cstate<=YUV_Nstate;
		end if;
	end process YUVCLOCK;
	---------------------------------------------------------------------------
	YUVmachine: process (Vsync, YUV_Cstate) -- clk pixels on 4th pixel, so they are stable for 4 pixel clks.
	begin			-- 02.07.07 changed Yclk, Uclk, Vclk, Y1clk etc below to correctly reflect pixel data order in stream from camera.
		case YUV_Cstate is
			when "000" =>
				YUV_Nstate <="001";
				YUVclk<= '0';
				Yclk<='0';
				Uclk<='0';
				Y1clk<='0';
				Vclk<='0';
			when "001" =>
				YUV_Nstate <="010";
				YUVclk<='1' ; --and Hsync;
				Yclk<='0';
				Uclk<='1';
				Y1clk<='0';
				Vclk<='0';
			when "010" =>
				YUV_Nstate <="011";
				YUVclk<='0';
				Yclk<='1';
				Uclk<='0';
				Y1clk<='0';
				Vclk<='0';
			when "011" =>
				YUV_Nstate <="100";
				YUVclk<='0';
				Yclk<='0';
				Uclk<='0';
				Y1clk<='0';
				Vclk<='1';
			when "100" =>
				YUV_Nstate <="001";
				YUVclk<='0';
				Yclk<='0';
				Uclk<='0';
				Y1clk<='1';
				Vclk<='0';
			when others =>
				Yclk<='0';
				Uclk<='0';
				Y1clk<='0';
				Vclk<='0';
				YUV_Nstate <="001";
				YUVclk<='0';
		end case;
	end process YUVmachine;
	---------------------------------------------------------------------------
	
	
END SyncProcessor_v1;